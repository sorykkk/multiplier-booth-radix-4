ENTITY tb_register_a IS
END ENTITY;

ARCHITECTURE sim OF tb_register_a IS

END ARCHITECTURE sim;